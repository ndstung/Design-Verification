package project273; //project273 package

import uvm_pkg::*; //necessary to include this package in user's package

//include all sv files

`include "seq_item.sv"
`include "complex_seq_item.sv"
`include "complex_seq_item_time.sv"
`include "complex_seq_item_fft.sv"
`include "complex_seq_item_fre.sv"
`include "seq_item_bit.sv"
`include "seq_fixed_point.sv"
`include "sequence1.sv"
`include "sequencer1.sv"

`include "driver1.sv"
`include "monitor1.sv"
`include "encoder1.sv"
`include "ifft.sv"
`include "fft.sv"
`include "decoder1.sv"
`include "scoreboard1.sv"
`include "agent1.sv"
`include "environment1.sv"
`include "test.sv"

endpackage : project273
